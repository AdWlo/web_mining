���      �sklearn.linear_model._logistic��LogisticRegression���)��}�(�penalty��l2��dual���tol�G?6��C-�C�G?�      �fit_intercept���intercept_scaling�K�class_weight�N�random_state�N�solver��lbfgs��max_iter�Kd�multi_class��auto��verbose�K �
warm_start���n_jobs�N�l1_ratio�N�feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�	responses��reading_time��publication�et�b�n_features_in_�K�classes_�hhK ��h��R�(KM��h$�i8�����R�(K�<�NNNJ����J����K t�b�B�                                                                  	       
                                                                                                                                                                  !       "       #       $       %       &       '       (       )       *       +       ,       -       .       /       0       1       2       3       4       5       6       7       8       9       :       ;       <       =       >       ?       @       A       B       C       D       E       F       G       H       I       J       K       L       M       N       O       P       Q       R       S       T       U       V       W       X       Y       Z       [       \       ]       ^       _       `       a       b       c       d       e       f       g       h       i       j       k       l       m       n       o       p       q       r       s       t       u       v       w       x       y       z       {       |       }       ~              �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �                                                              	      
                                                                                                                                     !      "      #      $      %      &      '      (      )      *      +      ,      -      .      /      0      1      2      3      4      5      6      7      8      9      :      <      =      >      ?      @      A      B      C      D      E      F      G      H      I      J      K      L      M      N      O      P      Q      R      S      T      U      V      W      X      Y      Z      [      \      ]      ^      _      `      a      b      c      d      e      f      g      h      i      j      k      l      n      o      p      q      r      s      t      u      v      w      x      y      z      {      |      }      ~            �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �                                                             	      
                                                                                                "      #      $      %      &      '      (      )      *      ,      -      1      3      5      6      7      8      9      :      ;      @      D      E      F      G      H      I      K      L      N      O      Q      R      S      U      W      X      Y      \      _      a      b      e      f      j      m      o      p      q      u      v      w      x      y      z      {      |      ~            �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �                               
                                                            !      #      $      %      '      (      )      *      ,      .      0      3      4      5      8      B      D      G      I      J      N      R      S      V      X      Y      ^      _      `      c      h      i      j      n      o      q      u      v      y      |      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      L      �            x      �      @      �            �      �      �      �      �      �      4      �      �      `	      �	      (
      �
      �
      T      �            �      �      H      �            <      �            h      �      �      \      �      $      �      |      D      �            p      �      8             �      X      �      @      �      �!      �"      �$      �%      t'      )      0*      $,      �-      @       N      p�      �t�b�n_iter_�hhK ��h��R�(KK��h$�i4�����R�(Kh8NNNJ����J����K t�b�Cd   �t�b�coef_�hhK ��h��R�(KMK��h$�f8�����R�(Kh8NNNJ����J����K t�b�B�J  ǋ,mrq�L>�u�5��@�~-��㿗��A^��z���(���DĤV&�?��b����B�Z�?3_	D��?0���. ��щ)!��?k�#��~�?F*ƴX������P�f?'ʭl6�?k"&��|��#���?�
���]�?��[H�q�y�����ĿX�O#:��?�.�t����x�V9��?��Gn�@�?D i�;��(�U�t?M�]?ɼ�?6����u��g@F@�W�?��lf���?b��?�� �Y��ծ�?���7�?��VZ�������?�q�#��?�&"8(C￬7_<O0�?Ce,��<�?�w?)��"hQCO�?O�����?|@%��9��IP���_�?)qjʏ�?�b}u������}I��?��4?�?,x��������|�?�o3,��?�/V��V忆�[cM�?D!'���?�0mT���8c
���?���$X�?��3��+��hz8o��?M����?������SE�e��?\��j��?H7K�́�qV�2�?d��rz4�?��7xf����w;���?�=��q�?ϊm�����C���K�? !�[���?Fo��3񿮎��?����J�?������+�?�!5�*�?1�|̐���H���?j�cͦ2�?��$�e�?�^У�?�V�Ne��?���o�]�(����?���B*v�?~�=�I��|�����?��_tU�?���{����f�\��?��mm��?��B�����_T�?v�z�XV�?��C��o�s�����?&�U�M��?8{|�R���f3h�ɤ������?)�.gw���
��?Zx�vI�?E:J]��࿞lO1� �?��dګJ�?�K�u��i��U8�?,�8$Vl�?�eR}O=�ړ@��`�?��y���?f�I?5�዇�i̻?枂x�?�oB��<꿂�2+��?"c��ޫ�?�<��%�mjp�c�?�1��p��?uR��A����.?����?�p@v�?��V����p���?>�D %_�?c�[<���k7��w�?8݊�`��?!oCH��ҿ���*&��9t� ���?|H>Fݿ�}�%#�?�d^U���?@�#�{���l��[�?�7'd��?�u��c>��!�E���?L��2�?UQ���H�3E��gM|?��&	�?0e\��ڴ��޹!R��?�u�E;��?~�Ţ�m����Y��?|��x���?�&��8�Q7�]��?3��Ζ��?B��K�N��,�?���Q�?��B����X���?��6,G��?���D���z|:{>��?� �P��?�֒(���d\��?cj
L�?\qPZS��X؆�?6�o���?�^�������(L�?5]9�?t�K�*��6�\���?g�'U���?e��6���>d��?F���5��?�W&���Avۉ�?.������?ܭ��w���S!�C���?y�.�	L�?�?/��x��CS�J�	�?-xC�_ѿ��ZU )�LP?Zm�?��S�@������xv濉��[��?4���$�?Rk��:�"���?M��k�?F�X�]�9{-gL~�?B_���?������ �G�>)�?7�m~9Op�� fː���^͈���?X��D0S�?Т�K����̃Y�ɉ�?��Phw�?L�O1����RN�[�?��Pe�?�?�~�W���P�&��?[X4g9�?�V��]�b��5C��?r��r�?�Uy"��'H\*��?�:"����?�#@_��!�=��?��C's�?Kxbu�ￖ�Yh��?��li�?�?hre���IJ�4�?�m�����?M����迷�z��H�?�&�P�K�?~S���󿻤>���?pM�ٌ�?������:��0�?���͠?)Y��ˢ��c����?d�����?�a�?��鿆�)�?�}�����?��)6wܿ�66�̤�?�m�����;	��2�?��9���?�K���F�^P��ҽ�?�~��}�?2���;p���O��L�?HOagc��?�A��T���W��?9U��^��?�L�#��Կ�K�λ��?6����S�?A���A���*���?&S  ,��?<�ޜ促Uc_��?���ͦ�?��_�W�L:�h\�?[�$�
)�?
���ٿ�"^����?�EF�~�?a�d�]߿�f#w2$�?��Ƹ��?C�-;���{�0�?��BF�?��t�ǭ�!�ݗ��?��X����?lYK%u��_'�W��?C���|�?4��`��㿤�r���?}pW�@8�?U F3������]�?0�$U��?N��������/�?���A��?vƵWX��rQ�Q��?�j
sݙ��L���T`���_3M�?ΨäK�?g~J��jB9��?\ LL��?�P2g׻忁�6xM��?�}X�U�?5 ���g�{�@tN�?�9�	T��?ȿ������#X�O�?�w��xk�?�q���(ݿ�f�?��c&��?�܇�(-���hmY/��?����? �h����}�e���?�z���?�@O�1�f.+���?�&�/vu�?��N�%P�ԟ-���?u�h��M�?�vk,|�߿^)M�s��?�q��Un�?n)����2n�e8�?:SfDY�?w�j
^�пa�I���?9]bWo�?������?te�(�?C�����?�[l)ڿv�R%��?U e0W��?-�R�Xܿ��wō�? g�]��?�O�y�ݿ?X'۰?Ti Sj��?O��俈 ����?'
�]�5�?�}�� ��v7|���?̯Y���?��lܨ���'�����;���?rqMz�׿�#t$��?�F���?���E��ٿ/n��-�?���w��?�CX'��¿UDsS}�?uq�%��?�J��,~���{��?��n�?e��v�c�GmOT�?-�]2l�?�Ӽ�+j���:��?�k���? �`㿌i�ו�?ʇ6����?	+4@���E<����"���?
Z̜V￸r��;&�?������?-�gZb������i�?O�I;x3�?�
�}�e������?&��B���?Ls�(��Ln"��)�?�����
�?�	Y�	�Pf�sDD�?��{���?z����L�28�/��?GS��g��?�@��cϿ��gY"��?{E��i��?AS��"���kC�4@�?u����?�9B��޿�����?���6���?v���ٿi�C�)��?���Eʥ�?r�L��Ŀł�����?��&y���?b;�rE�?fz�d
W�?$W�xҪ?6�Y��Ǭ�B�Fo[�?�s�p/d�?�����ҿ��]����?iw�,���?S���d�?����4��?��;X�u�?r����??�6�[�?�Q7�D&��F�7'U$�u8�?"�?2�w�?Mj��*տ�\���3�?i+�MD��?��, �����	���?vB��'�?+����ѿ�~�@��?~Z˜0¹�Z�h�ӿ%�v�l8�?3`�����?:
6���?�'��N�?�i�~!W�?O1ט�տ���_�?�x$����?6Y�3̿�j���?�IS\�?�w*�Yֿ��Y�? �^E��?m�<#}\п#�']��?����?p�e�����̗e!2�?&I��M�?��)چ�Կ�`����?�Mˬ��?�R���ҿN���`�?Ǔ�?��??�n���߿b�UB�?��<�j�?l�4���?TF6���?Pj*E�����"�3<�XRH���? �C��?�PC����� ����?:7R��3�?�G��{�ѿ���T{�?�7����?;^}'�?t�>Y7�?�#����?�6]�F�ѿ(ޡ�l��?��ŕ8��?*��و�Ҏ�<U�?L��?�T�肒���j��?4u�`��l?�z��3&[X�?����+m�?�u%4F�Ͽ����h�?Vw�ٗ��?l�#�k��<�rx<��?/��y���?�yy��п�ޯ� �?3��e�?{S���ѿ)P���o�?c��,4�?1I��EY迪H�����?���@O�?*c���?�~в����.#Ƥ�?���]տ���>3!�?N�°I��?��I���0��'!��?�c~��?^\��'̿鯾��xÿ�zO��?4�-)�>ɿq65o���?�}����?4����ӿ�P;��?��t@?�?J�q� �X�ƴ-:�?��ȬP2�?zx��}��@�s�zx?�������?ԑ"/��?�+sV"&�?rQ���d�?�>�����جj��?g�4]��?�N�L����^�Z�J�?��u���?b�-b�2��f1�!kL�?�Y�-��?&Y'y��?9A�(�?ӏ���?]����K��=�����?���N�?��MQ��߿�]������	 ���?�{�w�C��!Cf��?E}���?�	n��{���:�����?[Ҩ�Z���:��\��?����<F�?Oݰ*v�?��3ѳ�ӿ2E��n��?c�E��\�?�C�	*ǿ܆���O�?�f�����?2��ҿ�}�0��ɿ���h��?^!!D�ѿ����?�)��v-�?��r����?X�f�޿j�%��2�?}RL���ο0����?��C�_w�?q)J˜qӿ"���f�?6�g����?�����Ϳ����`��?)M9l:P�?'��f���(j"})�?{(O��u�?<~,��ؿ���!&�?5�����̿M��)����C�z���?�m��L�?7K��- �-�T���?/��a\�?�sA�y���s`�?�|�*'S�?��f�K�գx���쿔�����?�����b�?��+��?�ԣ��n�"��������ѧ�?
X�����?y:Ʈ���r%�^�?�z��L!�?6mІ�pֿ����*C�?}��6?j��.A�����o���?.�fV��?rr���޿�(A���~?Đ��?[٘[���{,[y�?ҙA7��?62�1wSӿݞ� S(���y�.:�?�S2���ο�
�C�_�?�5*$
��?I�d�������Y�Iʿ/(@^P�?c/�
R�̿huț�6ÿ+(��'��?0����]�?hO7Z1 �?�ǧkJ�?�/�w俿ņ�82�?��n���?ӣ��ih��R=T��?��'��?��MK�wӿfc�/I��?g��uN�?�b�iu�?����D�?��z���?r�9 �����{%ȿh��Z�?^��ۿ��_Ag�?�1����?U�t�6W��p9\��?��w�`����w����?��Of7��:U����?�]�Á��pN�hq�?���tA�?ͲYw�Ͽ�ES����o��+���?����OY�?�����?��;�.Ŀ����yſ j|����?1�ހ���?^�Z٦�?�1s�W��?��5r� �?�r�i�ÿےwTȀؿI��K��?�9�H����k�&�?������p5&dҚ?:f�rt�?+0Y�
����m��3⿑�1y�Q¿���M��?��t8��ɿ��N6(c�?d4����?�h�����?�.+�v��?@H݋H�ο1�8�i��?�����տ����1�?q�a�׿{����7+���?H�<nn�yn��(��?Q��C N�?�n�d:�¿S��>�?�#T^�,��{�$ſ;�UH"�?���y�?���<z�տY�z����?�gȳ|�?�|H�v�¿�!Tu)�?�>0�ʿ��A��ݿ��݌�&�?��S ���?�E�p4+�?!)oA��?���"�̿��B���?�^+�^�?�jj2���?��Z5��?ٌ��������k{R�?���@(㿲����?�2N�ҝ�?��8)\>��WЦ��ҿ߀��V�?K���'꿚���9�?B|���Ϳg���p����Yٶ?*d��{�?`���U^��a���X�����h�8�?8琀�Ɔ���J�?�*�����?�l3�`��?�L/�V��?�VD1�k��������?c6*���?���L$"�?�VA)�O���Ûm���?⼏r�?!3��?��;:w�[]�?���m/��?��~����{�����UH'y��?޶c�W��?
�	�޿�����?�.A�Tf�?{�<P�?| �R�㿓�A8	&�?����B)�?
UR�M�?˒���ݷ�8��/}~�?�_-l���?Nj��f��?���q�(�?+_�+j��?�<���]Կ�$,-��?��6n�GU����Ĝ9���ؕ �?w=��<������#J�?lE��-U�?mR0�"��l���?��V�)�Y�^'�?u��A�ɿP**!Pd�?�`u����?{��_¿�F�t�?-qa�&A���zYC���>G��KdʿW�\��|�?�0����V?��	c�?�U��O7��º�\{a�f�?��9Jx��?q����7�1��?�"����?Xq�m���?��V{��?<�&P���?���yS~�u�����?�<%0� пd����?�����?�=�ߙ
�?�%	�;��P<a<��?�	1�JJ�?9Ϊ+$ �?g��,t�Ͽ���m�����(���?��?ȟ0�?3A�����۳5l�?��"��?��*"�lӿ`ʬ?�����z>K�������?��9�+C�׼�=��?���7�1�?�d��S�ܿq�}C�?}K�)��?��r�i�ÿ��wTȀؿO��K��?�qn>fXҿ=,�`�D�?;���H�?r����?7��wϘ�?H�$_&p�s	k��"�HH��F�?W5�<��?2�p�U⿄�@Z�?��-���ڿB3���?ccè�����✻!�?�.0L4�?�kG&E�?"��6��?�T)@���� ��?�oDe[�?�4J���?�X},a,�?~b��q�?��h�3�?K3'��e�?M��@$¿���W�j�?�M�$�?���Xs�?����?����'�?�������:�˔<�?1��h���r��X�@�?}�T��$�c~T���dnp��?��/���3(A�?�O�P���?l�`IQ��+�'uӆ�?�r9 [.���E���i��z��?�T�� ��o0D�vp�?�?�� ���*	�{ס�?,G���?�_�fϿ��Q���?�/=v��?n�X"	��?k/1�c¿j.�b���@����1�? �x'���	��v�����Lυ�ѿ�d=�H7�?0�K�˿¿�G,�q��?�G�,׽?M�R�׿��h��o�?����B��?���g:��?�I��ÿĂ��ޔK��W`�q�?�<�|��?7��ˋ�?��.}/l�?.�xB�?Q���Ϛ㿴�v�]Ӕ?xi�����I_P��?�����?��i���??��d�ǵ�
d����?�[qb�i�?=�oc���x��LԻ˿���xj+�����yje�?��+��s����8�s�?����^��?/<��ӿ*!���?C��u�?% �]�?��=�{�?�[_y:����y�ȿ�?��8�ة���p2��?�S=[�8ѿ)sdRڛ��z����?7Ӭ���?�J]+9h���Ӎ�#��?������u��L{��? s�jt3?J��(�ÿ��9a���?�x�?M�?���%�ؿi�`��0�?�� c`��+/�rʿ�6����?f�	�s�?�n��	�?�h��
ǿ{2��&q�?�.�����?����E��?7`q�
p���S��+�?�����?:M�E�ɿ�ejɌ�?n@jt�?�����տkby�B��?�s/��h�������_ѿvv�PJ�?�"nh�s?���Z�=�?�� ��Xȿ���c��пUmL�r��?�X�M��ѿ0��tm�?*t�d���?�\�(k��?��CʯB��ajR�4ſy�}�7��?��_�e�ɿ��S�M�?(LK�r;�?E*N{d�?��V̿�Eh�bh����˼���??+{�8�?�4�P&��?���-�Cʿ	lg{�?p/*I��?~����y�?� EQ,ܿO��F��?�&����?��6�п���[�?L@����?�͹�忿�*~H8�?*h޸O�ٿ R�a���?z8�>�S�?-M"�]�?����@ݿna�_J��?&��˟߿ ��ڪ��?:���l��?��\��?[�Р����1��¿�Yj��2�?�Gv��ο?&tQka��(Հi��?C��SۿG�(���?�H�t���?ZC 4Oؿ4=-۲�?Ԋ�M�N�?0�R_p�?*gf��Ib�L~Y7Pn?�4h�A�?�)��?uH5��x��n�z�Fe�?ܡ�'9��?��(^��?H*יE��Ey ��?ȯ�Y�V�!q��	�?��A�q��?V':!��łc���?n�_a���?�HDؿ���ɱ.�?&�������"i#�?"�r_�?�b��J��o�0�B��?�ɇt���?P���?��y��?r}�U��Kjm�?.shՎ�?�^��׿��x�>�?�D�e�C�?Ĕ��h��?ώ��<�ٿ5
�����??��zC7�?������?劭��ο�s��h��?�b��:�Zq 0�s?,�e6%H�?�x+�7�?� �_� ��t+J��?C�v_/�?%;��?A!Z��9�,�b>���?J�!|����`����Ϳ(:���k�?x�-���$�+Z�?�Y�E�(�?���F���?L�IF��?	��v���
�Lυ�ѿ�d=�H7�?�R)M@t�{}����ɿ�Uz��?!7@��?�` �F�s�'���oc�?���.����q�K�?���Ņ�?ʲ�*J��?��ν�пx�]���?ŭr���ÿ	/&1x��?{�� ��?�}�jܿ��*�4�?nzT���?���W�?�'y]��ؿ��5���?b�h+���?�&>�>Ÿ?D1���?7�#����?X�B6c*ݿ|��{e(�?&�������
�q�u�?H���V	ǿ�!8G�lĿ�<��Ҙ��<0�����?���W�?�'y]��ؿ��5���?cf�K��?c�	(���?�G�җ�?𽅥6˿k\r;���?l�����uD^�?]῕�� a���5���?P׀Gf�?�M/�
&�?m/�;4�?���
�N�?�w�cٿ��Q�?m>�1wq�?�,\~��?�#'�+��yV��z�?Hbn�ȿˉ!CS��?��M�-]���s}�?���0~�?	Y{`�?���P�_Ŀ��w��J���\�(k��?��CʯB��ajR�4ſY?A	E]�?��R�?��J-{pȿ&�U���?�fSS����j��N�?�c��0X�?8������>?1KK�?t����?�8,�e8�?�C���?J��e�t�?�7���C���������?4��@'�?o݌ڨ�?D!��^濷�:�����U�?��pL�㠿1�>�t��?��	�]d�?�r@6s�ƿ}�T����c~T���dnp��?͓�S{�?sЁ,��?�n�9��?��uy���󌂜��?Qq��ʿ�������?��]�H�?#i�m}�gG
BR�?m���\(�?��.�*��xD^�?]ῠ�� a���5���?�U�E�?R�db-�?af��wÿϷ�R/��?EJj���?��/������S�����S���#��?ō�u�?h��I��?�@�����?w��_�?0P��̷����Xҿk�&欂�?T<��\��?����	D�?Z���3�[]&>>�?�d`�f�ƿ�"]
u�?���˭%Ŀ�~7B+B쿒�	ϵ�?�w!W���?��AXB�?"ؼ;�FпA���y�?��Y���?w�y�.V������俜��L��ǿ�����h�?��*40�?��'_&�ݿ K&�h��?_�ԫ���?Zj��?�����Kٿ�%@���տ�B�B�<�?}��#>K�����b�?��� �?���[��ѿ[%j���?��-��ٿ�I��Q�?�����I�?��c-�?e�~�Q濆�=C�L㿕��hn3�?u_�3KN�\�+32�?�����?!w��Kѡ�{�	f�ȿ|�r�m�?����A�?݋Q�D�Ͽ�i���ʿGNޟ��?�A����?Y2��Ȅ<L���?��*~H8�?Ph޸O�ٿDR�a���?N�� =\�?4.鰙.�?�ړOпQ���T��?��	�hҿDZ�����?S��5�C�?�d	`�]տ��$7��?������?��J[r��?k��ͬ���r���L�?e9(��'�?��$}���2���&�?��"bK���v�ݞ8�ǿ��,^��?��Mfƿ����x�?L漒��?�8�E]����9Ĝ�?��9��Q�?��؄ÿ������?�[
�?:�v߀��?��YFC��t5��?�c�mv���hl[!#p�� ��E�?�čt`�ſ=bء2�?����`��?�������?���8�[��<^ 5��?��LG\�ҿ")MQ�h������3�ؿZ��x}N�?K����?�o�4���@�>��?��6� ��?/�D�m)�?�B�!��?�� }	ѿ+i�H���V��7�o�?��i�%�ӿzi�[���x�K y��?7������?�����ۿ�莾�z�?���QK��-���̎�?��Z i�?I�ia�? Is�?�l���뿚��6�P�?��(Χ�?�th.�V��	��Lٿb�Th��?#�&���ſ$�wl���??T�a��?�^�g�?]S>R�U�?Sa�O$�;�t��&�?3Թo��?Ӭ3�?���J�hÿ_(^ӱ�?x%j���?,��-��ٿ�I��Q�?��4X��?���R���Є��o��?}���)��?��T�����7���?E�0'�&ٿ(1�p�{�o�QOQϿ�=[�?HE�N� �~Q�?fn�h@F�?tL�rտ�Y:Ns��?y����?/��wϘ�?B�$_&p�[��:�ܿ���`��?T��U��Y�%XH|¿ӫ޸��?����u�ο�Bc)c��skֿ2����c�?�Aq ���?��}�Y�߿]�����?@���?J�7s?����Z 6�?,�4��B�?b����9Ͽu��G�տ���a∺�zP�Rsp��]���Z���gk�n�?u����?UR�1����~6�Z߿lrY�
T߿�f��%��?y	��#�?�\E�9'�?�s{(+ٮ?̏���:�'`�*|#�?,��4xJͿ����?._ �(ɿ�p^���ѿ��`��?�������?���8�[�����a∺��O�Rsp������Z����UF]�?NgF>r�?EO�Z��׿����)K�?L�{6�ῈK��q�?�{�)�9�?�~f�3�?u&�ϡ�ￃ�8*��?4N�%ֿ�l�[���?��r�޿nR�h����(a��?�u�e?��?ɇ9�-�?O05� ����m7��Q�?$�4[T�?2���w�v�8ߒ>�B.o͋��?n�y�}�?�u��D��?��c�̙�?~�ȅ	ſ�-GWsݿb�ġ��?�F�G�9ҿ�~�	{�?7#�I���I���?ir�U��~���K��?M,��W3�?^+3"�
�?ļN"�����'h�UQ̿\�\uV:�?���n��?�iZ��eѿ�v6��}�?�OM�&ӿ��t^FN���9�K9�?(���f�?�m�gпnk��եؿ���d�?|O��p�?Rh!D:wпT�c���?A/F:�ٿH#) i�?�1�q���?��wuaؿ�z�#�?�R�慄ۿ��v��ʿ�aN9J��?@�SL���?N�$�/]?��(���*9P���?�����Կ_��ݞ,߿�w��Q�?qX��J�?��Eϓ�?pHH!��˿V�]QH�?V���Yf�?��@E��?�����ֳ�ؿ�#���?1F[��ۿ�D���?�;�=f1ѿ�w�L�ɿI@��d[�?A��8��?�I�a���?�#�����d49ӿ�Go	Hؿ�;�C�?����ά�?��C��W�bs�o�?!�{�7�?Wqk`��;?���T�MX��?f�����?�g�A��ݿ+�]Dh�?�~7+�?�-5����?���?7�D�?q/�{��ҿ��j3中��Y+�Fɿ�����H�?#�"
|��?��"ݖ<Կ���7f㿷�Y���?nU�8���?<�0��ʿR�@�hĿ��(ձ�?�x�w �ۿ%�;�t�?Pd�L���,�B2�?��ŒN��? �܁A�?�=L7�=��6�����2�_������Uҿ���{,��?5�
U��?����;�T����u�G/����?�j ���ֿ��#�_<�?��8Ui��?O#���ڿ�l �,ѿ�ݵ�Ҭ�? lP���?V��ٰ�?z{��F˿��+c�i�?�cD��?V)X~E�?q���L��o$�Vs��?��M^��?�����濥��rU��?LhX�k���06r�י?M��Ƕ��?D����տLHJNC��I��OL���D{cվ�ƿ{�In*�?e訦�$�?HB�R��?<Z;��"ÿ�v#%��?Թ�����? #D�4׿:�)�̮���1 ��ͬ�=�)�?���;�?�����sؿ�&���>ݿ �)���?�t��m-�����1ݿM�oi���?���|���?\�o� ƿ<f�$�?��bS��?��*��n�ދ�E�?^čt`�ſ2bء2�?LrB�ӽ?�a*�Iy��d��^�?"p�1e�?tQHJ&��?.4c��ӿck����?$F����?rT���忀p���6�?c&���B�? �R�ѿ�z�#�?�R�慄ۿ��v��ʿP��\��?�u�d�����7[��߿3������?�e��dп@S�}���?�/d�t�?~����;�?N=�.ٿ*NʽS1ڿu�aQ�y�?m��<&�/�5ә�����P`���r+K�?#�iG}�?�9nx�p�?U3"�ʿ�8�/���?��B���?����	hӿ��ɭ��?�0My��������?��9;�?��8���Ͽ�w�Yի?>�#����?i�B6c*ݿ���{e(�?2]Un��?k�Ye�����n���p�?e�_uԿ1V�$���R�h�]�?��q4�'�?�2Q���?cI���뿭c��pÿ�Y����?Z�5$�ܿ?�nJh��?�Jf�h��?f����wjH/�\�?�� Oѿ�I��v,�?���YH�?WE�[^?׿��z��?��[;:�??�ޝ���?M�y�8z|%��?"}�r ˱?v7E8r2�?�U¬[
Ϳ%��� h�?WU���޿�L2�޿F�G��i忁y����?yjH/�\�?� Oѿ�I��v,�?�0.�f忓]�oָ�G���Y�?�G�O)�������?%���%ݿ��j3中��Y+�Fɿ7����H�?�7��ޒ�?�DlG뿊�WÜt�?�׃lB�?�P7Ŀ����D�?�\�(k��?�CʯB���`jR�4ſQ���?ꖟu���?�эI��Bc)c�P�skֿ�����c�?+3"�
�?ļN"����\'h�UQ̿��"���?~c.����?�'n@aaпi~ S��?��_N�ǿ�ُ�u��?-���-��?tͨ����?��B7�ֿ���`��?�������?ɯ�8�[��h z�\׿��ѧ�2㿞��9��?P��\��?�u�d�����7[��߿�d�� ��?M��G�?�(e�������E�?D�����?DZv@"ۿ�XhDb&ֿ�#f?���? �������+���إ|m/���l;���?�+*��?iF�h�?bn��*���aN9J��?E�SL���?��$�/]?�,[R�?t���
�Կ���dۿ�k��եؿ÷�d�?�O��p�?�E~@w�?e�Jp��?�6���G+3"�
�?ܼN"�����'h�UQ̿�jwp��?���Ld�2�^|pv��u&���?cs��MJ�?4 c- �ӿPNq��vȿ���+%~ӿ#)�o�[�?�m\���?6�w�>�xݰ[�?D��9}=�?I����߿煿nfoѿ�l�����?ѭ#L� �?�\{����4�6����?��Ap1տ�keo���s�w���?�3|�?2�.�V�e��ІI#��?��%�X?w�����!N�[*��?�S�1*���¬]�?@��)��?we_nk��?�������Fa��?�c'p )忤���&��?|^#�ʆѿ�G��gѿ��}��4�?��ɇ-�?lm�]wſN��X��Ŀ�0.�f忰]�oָ�	G���Y�?!
�p'-�?ƏX�z�ٿ��T�ƫ�?��w���?�S^g��ſ����¿3��R�? �W� 0�?��}Tp�#(F}_�?��>f鿿7�8��?Y&J�Q5ɿ��Y82��l)NAh�?Y�_��?���Q�)$�C�|ֿ�u&���?>s��MJ�? c- �ӿ�l �,ѿ�ݵ�Ҭ�?�lP���?T+3"�
�?��N"�����'h�UQ̿Yl܌;ӿ5(���+�?��p�Lx�q���O�� D�jB뿟��b�?%�0}�? �D���?��R����95�?�Ҹؤ��?�t�Ìǿ�v�_�?]W8�G��?�oZ諨ٿ�N���?mG����ÿʟK�D�?3+3"�
�?ȼN"�����'h�UQ̿�i�����?0#M2��0z�-��?-�4��B�?.����9Ͽt��G�տ.\$Y~ż?!�N%�ه?��m��ۿ��9�+C�м�=��?��7�1�?ø��G�?4�
3�����smR�׿TDW��5�?�}����?�����=[�?"E�N࿪�~Q�?#�4��B�?����9ϿB��G�տIf�$�?��bS��?��*��n��t5��?�a�mv���gl[!#p���Fbơ�?`�F�+���@�PV�ſ��Ŷ[
�?���2BR�?{vMm!��F�W��?�B��#zٿ!&+F�޹?@���f/�?[M+K��Ŀ�s=����?]�%XH|¿�޸��?����u�οb���H�?��]�?^��q��=&J�Q5ɿ��Y82��l)NAh�?$.QJG8�?��~ޯ�K>@X�\��J�꒱ֿ!}�?�?{D9�_�
�ʄG���OϿ��-��?1a/��?��!�ÿ׿<.�_$��J�v�yC�?�k�y�Q�?�SXқ���E-P���?���Ա�ӿ�w�zIB�?F0f!gT�?S_�d@�?v�3�6s���i���?���X�Z�2L^W๿!����?�	��ѿ�˥E��j���G�?��S�q����~hjSu��G-��N�?�%�p��k�]�z���ܿ��#L�?.�R��?�;/�Kh�Sa�O$�Z�t��&�?:Թo��?<�u�c�?~��A�?'p>˲��;��?*�?q��Y0ٿ�	����ٿ�,[R�?V���
�Կȵ�dۿ:0%�.��y�wk��?E�%M5�ʿ�z�#�?�R�慄ۿ��v��ʿ"�ly\�?6B��]���ޣ��E�?�0�� �?2��#�Z�����+��U#<yXe�?���)Q�ȿ �3�iA�?�z�#�?�R�慄ۿ�v��ʿCM�9�@�${�:��?�����忩r�p���?���R���?1��p��¿Y%j���?5��-��ٿ�I��Q�?iyT8�W�?��la���=�:5���s�nH��?3��1�?���um쿻h��e,�?���J�¿�������/d�t�?_����;�?,=�.ٿ�B�Q�m�?R�0�D��?��?���� ��B��?�	\ک�?��)} #������t�?��j<���?�Q��|���he���?���W�?L橦�bȿ�@LZ]��?+�!e��?�vVG����eK�T5�?�a����?0(	:�t<}O��?0��<h�?$Jq�D�4�~� �?��\��T�3��{:�?��JU�?�:a���?up���ɿUa/��?�!�ÿ׿Z.�_$���?P_��?�� �>��L�s�Lrտ
�p'-�?��X�z�ٿ{�T�ƫ�?��F.��?TJQ�$�?+!}�C��ڋ�E�?�čt`�ſ;bء2�?6^ 5��?��LG\�ҿ�)MQ�h�������?�+��������])w:տ������?�����?����ճڿ�9N���?c迤@�?��k �㿜%@���տ�B�B�<�?��#>K����o��?�Ut�2ֿ���d�?pAQ�翦$Q���?kl�A�������>�?4J��DJ��%RX��?�H�NG�?N�=�&̉��"W�j�ҿ�:�[�S�?��c����?߈�RY��A�=���?r�P���gk.i�l�?ǲ?�5�?J�gU�¿5�S%�?ěu���ֿ�˔��*���-춮��?0��*��}?��W{>�?�TK��ؿ��%F��Z�k �?����[���~� ο����9�ܿ�W���?̏���:�.`�*|#�?��4xJͿ!�J6��?�?�q9٬�ަo𿫩�a∺�hP�Rsp��z���Z����.�\;��?v�)���?�O�1$	ݿO�,���?T
�xA�?�+��տ��$!=��?�Ks�տ�����W�?r���6��r�"ɡ�?�9���ո���#��?Ʋ��5W�?��q��yܿ갉�x�ӿ��P��?�)��l��X��C4�?Q���?Կ.)�ټ�ٿS'�
�z�?���/��JW�0�𿷜�	�?�h9��翝C��?]|rK���?��&`���J��@�خ?�)�֥�?���`[�?"��:���6� �c�?�$�Z~��*�j�	����c>dU�?z V�����
;��Z�̤�ۿm_-@p�ÿ����v�?]��|T��?3�!�X����Bs�ܿ��bs�5�?�b�3���?{BPG��fdw���?�'q�	���u��L����^��?k|���(ҿ�󽭜�׿`�	's�?�����ȿ>���!=����v����Lυ�ѿ�d=�H7�?��f\��?���W��?Op����Ϋ��?�	��ZJ��}<⤿�7��ޒ�?(�DlG�ؗWÜt�?�e��2$�?4�s����?.^��=�ֿY���Xz�?gT�̑�ڿ��n+kg?��'(��?Z�a�G���ݟ�f�?���ۍ]?k�Xx8b�?�r�ֿ�n4$�"�?����w�?fe�[,����i���?{��X�Z�jM^W๿b1�n��?���.?п 6��w���TQo�S��?�
Nٿ-�ް��ݿ���^��?w|���(ҿ�󽭜�׿ɲ5h�2�?Ve`�l��㭭<�ɿ���g�?8#�;����>�}���n#c{�?�^t:{�@�$]A<�?�~��lb�?�X�T���?`nS'~��|rh�Ƕ�?��`�A��?d��P�Կ��Vw���?8I�ш�?�Eh�;�?�Ry�H��?y�!5�O�?�#���¿p� G�B�?�^gQX���)V���ؿ#���?r������?o }p+�׿�w>|�?����B�?S����x���K����?Jsrת�?�-|�E�⿁$�b�[�?z�Y�j��?n��<W⿠�-
��?���i��?
��W�L�/��!���?)z'"/(տz<���ӿ�0�� �?!��#�Z�����+��z4˂���?�%O���?ԍD:���P��K���?� @��wԿ?MK�7ؿ���l�)�?�J�ٿ�)��Rpտ���X	��?2aY?�?�B��ҋڿ�����?A�\��?!�w�M�ӿc�M���?�Xu�9��?��Mc\޿�@�\L�?eY��Z�Կ6� Z�:�?������?G־ �B�?����s4�	��A^�?r��C:��?��(ʤ)鿫���G�?y�_�O�?���G�Կ{�F���?"�F|Ǩ�?s	)�)�Կ��\K���?�*����?PX�Y뿳a�/�?�|2��?D�tՊ#�+��9}=�?=����߿��nfoѿ��m5-��?����G��?�����C��B|K�m�?��_���Y\����㿳�!K��?s�Y%�Կ����>�A~W���?ڋZ&�c��Gq���tÿj��3��?���i��?P�ݡ2�ڿ8�/�i�?U�<��?O�BT��`��y�?�����n�^$������6m�?���/ވ�z@)�7�?#�$���?��q���?"Sx��d���� �^�?⸊{}]p�F�����ֿ(���P~�?O
�
��׿"��.Ͽ� ��?������忆M�5-z�.FùT�?<^�?��?��OB��i��٥�?<���u�ҿ�XH��*���f�?5\h#ٿ��s
g�����G��?�P(f1����ٳh𿔃�Kų�?�*"v�X�?�������kh����?^�ۿ����C��K�rW��?�C�w���B�|��c�<�S�?U�[�2�¿�o���7.�����?U�]�����ދ�� ���$J�?�?���6~Ͽd���|�{����
h2�?�~�zo￷0����+�,S|�?���4��?���������8�S�?-���K��?�Gܠ*K ���M��=�?��`�6�ܿ��p�/忲K��b�?+.����hcp|qiݿK�C��?f�f��?�&%���غ���?u'R🄿����濋گ�|j�?�HL����J�㿉����?'��ܿm���)�?<�����?χ��Z���<Z�_ܿ�)�?}��?�P&��ۿ�6��Jm���ѱ� �?2��0@�c�8-����4|�J��?�"��z����,��?b!�Ye�?֪Z�����Վ+���i���?ܪt�������]��鿱��3��?�c1{M��SGό���E~�O��?z~P\������d�nD�"�z/w��?�zi��~̢����_H����?���Ǘ.��D�� �t�b�
intercept_�hhK ��h��R�(KM��hN�B�  H� K@	E��`@Cy�0i�?�Ҭ^@��?:Pl���?j���L�?�[Ā�_�?N@]��c�?���GIǿl9u�{�?�����?(�^�֌�?sl_�?�K��S��?Y�&���?�廈�{ÿ*������?s�p[MV�?=�V��?��m�Ց�?�hnn�-�?�c`�L��?�\co�?	AW1X�ؿ���V�?��(�#^�?Ε�Yv%�?�QN����?+]Իc
�?�-�#1��?��Z����?w>KS��?�񝑢z�?o�TB��?�w!��
�?�ΐ�w��?Z�?��t�?S����T�?�Vb��缿_�%��ؿ���t7�?�Nlu�?]{/�!��?����T�?,OlJ���?�Q��6#ݿ���B���?y&7���P��i�?�#����?A*{?���?�:�v@U	@��A*4�?�3�T@Q�6�g@�d��"@��/����?�'�QT�?�� ��?�]'y��?�&�%���?_ۑg8�?;��)�!@!��q��@�d}N�?J*8	��?3�n�c�?}�]@3v��K�?���H��¿�	�R�#�?(�����?�؍�\�?WZ?G���?�W�����?������?嚓;��?�9ۯN��?Ӗ}ۆ�?g÷���?gW���?x@-��p�?��8��@1�/�y��?^Б��g�?�,0i���? mЬ��?��k��/�?�{r�Y�?UY����?�d-�?�c����?���<��?�Lc���?Ʉ����?X���׾K?�J�g��?�1�ZW��4�E��ݿ�2.M�?O�3�@p��1�?�N廭w�?�b����?����?G�*�G��?�tx�	��?�����2�?��b��?�o��i�?D�d�ȳ�?N��j���?u��^���?!qz�����r0�꿝M��_�?�e2S�ɿla1���?�v����?�ʌ6��?����F�?}����?�º)&X�?I�L��{�ؼ��Ι�?ɩ�$g��?|�8^E��?�$Q�f�?f�܆R��<�4�kڿ�0:���?R|R0;�?*���(d�?�=�����?xW�6�@�?��J�Gp�����m�9�?�B�b��?2�d����?Z����ǿ"D��w��?�Ur�G¿�������i�	�����S�̿$Wgk���Q�+����?P>��T�?�X���+����xr�|�?������?�\t��?0�i%�?���	 ��?��/���?ś�'�k�?�iP9?�??MnZ��?��|�s��?;V��ݿ�@q�?0M
�X����i�몿Fށ1A�?5��G�f�?d�ĕ4;�?�l*i�俏����?���2G^�?��n�f�?�i�j3�ѿA-�6L6�?S�V�P��?�aY�wfͿ6��.�?ɨZ'ҿ�z+g��?��K4��?�ED�?}��׿񨐊ge�?Gd�����?�转`2�+�=�G��<�`t�咆ſ��'�Ԣ��t�y���
A]o�'���U��,D���ȟ�G�Ϳ����ۿS~�^2�?�
P���e|��Cӿf.a�qeǿ9��g��?�G�'�L���0�?��2xִ�?x���R��f��
�����׽п�PZ|z���V����?����}�?����R�?�$���?���1���?n�DvKrÿl}�r�f�?v�}�?3�	��߿�z����?ѥ'j�鱿��t�t�?ϴ:2�ֿ��zj&�?�ۢ���;�؜�%տ�������?4���m7ſ�y��@�п�[{-�k��R�ai�IĿ�:1�"z�?�`;����?T�3?��? ��Pl�?����&7�?��j��?��u�l��?���m`�̿�$��{翯�<��?�L���d��N�z���?��~O1�����8��ҿ}����m��ӿ�y�3(k�?*E�G4ݿ0U���?�(����k�o��Oƿ��A���)pP�=X¿t�5��ǿ�S��4-׿�Qk�
ſ� Y��ϿZ�����F��+ѿŰ� �ѿ�+|�uKɿ	v� �ӿ=i�.b�?��z~kڿ�s:�@�忪�1J���o�x�"�ͿsOu������d}��?���?q��{�ӿڱeAJֿ'�H?��??ZJ�s1׿���;��տI�ɗ���?CCJ�տDhDD\ۿ���Qƿ�A^,��̿�4#�\������A.�?�W���Gο���[|�?�:����?�JB;��ӿ^1k�c�㿻���&7�?���7����&�g߶���&�_����#̿.;5������<�{$��?ܚ��2�?U�c��¿BYH�~¿��l���Ԓ�c�g�?�j�9Mֿ9�R2�ǿ��3��s�?j'�O��?k��C�,ڿ�t����?k����չ�ʡ��Ifӿ�-Y�B�BS�|4�����q��ڿe�8�V�ֿ��h�̬��W'3X���0�xz#ʿ�+Y_"˿��x��?S�fQ"�?�v �˿U�k�̿v]sAǿ��38��:yb(�տ{�ǯ1�ܿW�@���˿.5^M�ɿ�Q���Ͽ@o�
gϱ?�i>��c�/��oTG��N�.�;�?���m��?�ç*��?�GԽp����A�߳�T�Cq����� )d� ǿg��Ah��Jf��4�?�Aq��˿YDR�o�ѿ���ͳ���V!��?�5
�G޿�w��s�?�.�nr���n�g�8�̿}���@�Ϳ�2��^1�?vv����ٿB�S�?v�Zn�ܿE?�{�߿/E��p���=9S�?1�OlI[?��u�t��?��[4輿���И���PX��ҿT�S2x濔��&�@�?�JHk��`8�A�ӿo�3d���?��$�a��{�XG���������~��؊��!�i�)?�T�;ѿ$e�i�(ſS�|4����?�쯿+T�p���?ř��uÿ7��l��?��vAx� ��&�����9k�S��ɺ-�~m��k����ǿg��eۿ�W��H﷿"�9k�S��g���z�ҿ�G,c#ſ��_���%�6�����8�{�?t��=AM޿ze����Կ��'!�ƿr��/�&���f��Ah��$%=U�ſXu��п��A�L�?��L�qޱ�m.X� �ٿ�(�����?U�j�!⿸��i��ҿ"�R2�ǿ_D��C�?[���!�ܿ�>��S���`��v߿�_���C��/ſ(�k(I�¿rr�7׿1Hd��ؿ�8� ��п� �*g࿑�v�E�ȿ�A� �!��5�[�r�ۿ�Pטѿ^���E�?�b������T��+���^��c�׿�>N�=P�?(ц(�?����z��m�>A^N\ʿ�v�x�6ӿ�b[�Y�;f�w��A?�QG��Կ20�nr�����g������}�d���|r�Dcſ�2&�dݿK�m�8����nQm|�ؿq
���?������?����eؿ�Z����ؿ���}�ֿzG
Efʿ��J�#Ϳ�c��u�?� �!ܿ�M��wOۿ��s"W�޿ո������f3� �	'��b�o�}�Y���͑�轠n�P��V	Jl��?�=�E���6
�Ͽ7�ޟz�?�ц(�?����V3ٿ�ϕr��?m�=�pɸ?wm~g�/ɿ���H�ÿ��&�g߶�9�������Z�yݶ�N�9"�M�?� ?�ʿ��ak�ʿ��b��K�� �Zi���f��8��=^&�����E���b߿�<�������J�#Ϳ�Zi�����~K��ȿ�,j��6ҿgRq��]�߷�ÿ>�,y�������ܿ�f%p����+���տI㲪�̿�KY���w��3s���П�8~߿�D��)�IV������*hI�?gX����׿Y��nn�Կ�4&�2mȿ���������IFe����˒�п�7�6�����x������P�"7�?"M%���޿]9�*�οq�:<�?B�ռᵿ�"I��ɿd}�!xۿ�-�Z��ƙ%X�w�����OԿ*��qҿ�E��<�?8�E�Ͽ5;U��7ֿuB@5[
㿋I�竹����Z2#�?�h��l�?�����d'�%b��?ۀG�ѿ����Pп��|�տ��D'ֿ�.��d����-�Nc�ڿ���-p������lɿ�ǝރ׿������῍�T&���?0ٖ�J�Ŀj�s��V�?�N��C(}6��ȿ~G
Efʿ��!;��ÿ��8���ݿGb �^��7D8U��f��IFe�����i��ſ�愄;���}N*���!�oB�?��Ĳ�ڿ���/#�{6��'Կ�o�����PX�?Q����ǿ.�/�s�ĿJ��rEԿ���ŕ/ȿ�!���߿�t n.̿ <-����ީ5��ѿ2��A�Pпhq���uڿ�uɸ��ʿ�m�O� ���;-����=����ӿ�1��ޞ���E��<�?o7��}�ɿw�<uP,ڿig��Ah���F2�Ńſ��9"�M�?��D���2��$�ݿ��W�ڿ�Sm��~����J�#Ϳ��T3 �տ���i��ſXIYX�ݿ�E�V࿷Ol"Qؿ.��6K�?x̩�N�ҿ���˒�п�!�ฤ��v��nn�ԿI~9b�X��S�D��DJ� ��?	�3�.v޿��vs���F����?Dj4wư�`n�H)��?SyG���H������%%V�?ԗ ��k�?rK��1S��\g�����z �]Bпy���'�?[����ӿܱ�ی�Ŀ����LL�?����a1տM.|_��ӿ��S�IE¿Ɗ=>����3�.v޿����Pп��D������
�NL|�ߴ�E9vj�ڿi��Ͼ�տL�|�>�Ŀ=C�t��?��D���HG�ϲ�?h�b��K�����;s��?KB;��ӿSg#W�޿�L�(wԿ�m~g�/ɿ��b��K�� (}6��ȿH��}�ֿ��*�`�ɿ�"�����n�@n�ӿ�2�ؖǿtZ�yݶ���v �ӿP�S�IE¿�iU�V����v��?l��=�Ͽ�|�t�g¿���"�տ�I�傡�OK4�ֿZ֑�y?d�О�]?HN��Ϳ#C�p �տXR $�ҿ�6
�Ͽ�>Ĳ�l�?�$6H�࿾!�ฤ��4
M������IFe����YZ	ѿm�����ο����ƿx��IFe��%Ay}�Կ"���#�ٿ�І(�?���8���>⿎B�6Ď�?�U5�ǿ�N*�����\�I���q��GlտB�͉�࿻�{4�׿�#~P�~�?-@0�����w��ؿ��.	Ϳ@�c�O�ڿ�|�t�g¿� �r�����ی�ĿnWXM&\ܿHG
Efʿ2c��u�?35��˿���חῴh-��修^��c�׿�꫕�Ŀ�~������L�����{ ��ɿ6��V?Ϳrn�[�?�|����ſ��1E�ؿ �{
aĿg�\F�׿2A��8ɿM�b߿C/!���L�Zi���@�utL�ƿP!H����u�ѿ�D�WٿF�-��������o�Կ�<.啺���$�}�	���b�:|ҿW?8;Mh����D�Cῇ�c�k8�?8�y*?a��P\���K�?�R���ÿ�F�A�쿮��6�Ͽ�NV;�����H�(ԿbS�|4���:���l�����1`�?7��}�ɿ��V#)ѿ���aӿ��D"s�Ͽg�}�mտ���翩�Y֑�y?���	��?���.ſ�NV;���_�K�ө���v�[��g��֥�H?��'s��ؿ����?�up���ޛ�J.�?�hv���?��3��?�SVOֿ�s�Y�� �q�ܿ�?���?a�x7�B��������ο�!)�ٿ'8�x/�z?�eP��ҿ�(qa��c	���߿@�fr:zڿJ�|U�����u�<�L�׷j��� ��S�К71�C�RLc���_kK��j4wư�� :u�꿇��R�>ɿ\y)���f���(����y�^4/
#G�w!l� ׿_7Ua<Կ>�ᱥ��T���i޿�V/�X�ſl�8�N�ٿ�$�)@ۿ���b
ֿ��l�*�˿�}���[���n��q.����ѿT�W�Z�޿�	e����܏��tݿ~���D޿�5�v31޿o�S4 ��N``���]ǚa��ѿ=#3�Eƿ�2p1�俥1;C�:�5��xͿߛm��ۿf&h%�忀kW4���z������y>iDܿ	�IĿ"#x�x
׿�k��q�ԿMVdRcѿc�%õ�ڿ�Z��H^࿔t�b�_sklearn_version��1.0.1�ub.